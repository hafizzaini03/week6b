module seg7dec (x, y);
input [3:0] x;
output [6:0] y;

assign y=
	(x == 4'd0) ? 7'b1000000:
	(x == 4'd1) ? 7'b1111001:
	(x == 4'd2) ? 7'b0100100:
	(x == 4'd3) ? 7'b0110000:
	(x == 4'd4) ? 7'b0011001:
	(x == 4'd5) ? 7'b0010010:
	(x == 4'd6) ? 7'b0000010:
	(x == 4'd7) ? 7'b1111000:
	(x == 4'd8) ? 7'b0000000:
	(x == 4'd9) ? 7'b0010000:
					7'b1111111;

endmodule
