module counter_4bit(clk, reset, Q);
input reset, clk;
output reg [3:0] Q;

always @(posedge clk or negedge reset)begin
	if (!reset)
		Q <= 4'b0000;
	else
	Q <= Q + 1;
end

endmodule
